

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.display.all;
ENTITY DOOR_TB IS 
END DOOR_TB;



ARCHITECTURE LOGIC OF DOOR_TB IS

SIGNAL SWITCH   :   std_logic_vector(5 downto 0);
SIGNAL TRY,CLK  :  STD_LOGIC;
SIGNAL LEDs     : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL SEGS     : SEVEN_SEGMENT(0 TO 3);
SIGNAL UNLCK    :  STD_LOGIC;

BEGIN
DOOR_ELEM: ENTITY WORK.DOOR(BEHAVIOURAL) 
PORT MAP(SWITCH => SWITCH,TRY => TRY,CLK=>CLK,LEDs => LEDs,SEGS=>SEGS,UNLCK=>UNLCK);


PROCESS
BEGIN
SWITCH <= "000000"; TRY<= '0'; WAIT FOR 10E6 NS;
SWITCH <= "111111"; TRY<= '1'; WAIT FOR 10E6 NS;
WAIT;
END PROCESS;
END LOGIC;